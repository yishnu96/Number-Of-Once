----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:22:14 11/15/2018 
-- Design Name: 
-- Module Name:    SDF - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SDF is
    Port ( I : in  STD_LOGIC;
           O : out  STD_LOGIC_VECTOR (3 downto 0));
end SDF;

architecture Behavioral of SDF is

begin

process (a)
begin
case a is
when "1" => O <= "0001";
when "2" => O <= "0001";
end Behavioral;

